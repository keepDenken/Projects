library verilog;
use verilog.vl_types.all;
entity pr1_vlg_vec_tst is
end pr1_vlg_vec_tst;
