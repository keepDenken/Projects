library verilog;
use verilog.vl_types.all;
entity Project12_vlg_vec_tst is
end Project12_vlg_vec_tst;
