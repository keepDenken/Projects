
module mem32(clk, mem_read, mem_write, address, data_in, data_out);
	input clk, mem_read, mem_write;
	input [63:0] address, data_in;
	output [63:0] data_out;
	reg [63:0] data_out;

	parameter BASE_ADDRESS = 52'd0; // address that applies to this memory - change if desired

	reg [63:0] mem_array [0:63];
	wire [9:0] mem_offset;
	wire address_select;

	assign mem_offset = address[12:3];  // drop 3 LSBs to get doubleword offset
	assign address_select = (address[63:13] == BASE_ADDRESS);  // address decoding

	always @(mem_read or address_select or mem_offset or mem_array[mem_offset])
	begin
		if (mem_read == 1'b1 && address_select == 1'b1)
		begin
			if ((address % 8) != 0)
				$display($time, " rom32 error: unaligned address %d", address);
			data_out = mem_array[mem_offset];
			$display($time, " reading data: Mem[%h] => %h", address, data_out);
		end
		else data_out = 64'hxxxxxxxxxxxxxxxx;
	end

	// for WRITE operations
	always @(posedge clk)
	begin
		if (mem_write == 1'b1 && address_select == 1'b1)
		begin
		$display($time, " writing data: Mem[%h] <= %h", address,data_in);
		mem_array[mem_offset] <= data_in;
		end
	end

	// initialize with some arbitrary values
	integer i;
	initial
	begin
		for (i=0; i<7; i=i+1) mem_array[i] = i;
	end
endmodule
