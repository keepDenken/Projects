module control_single(opcode, ALUSrc, MemtoReg, RegWrite, MemRead, MemWrite, Branch, ALUOp);
	input [6:0] opcode;
	output ALUSrc, MemtoReg, RegWrite, MemRead, MemWrite, Branch;
	output [1:0] ALUOp;
	reg ALUSrc, MemtoReg, RegWrite, MemRead, MemWrite, Branch;
	reg [1:0] ALUOp;

	parameter R_FORMAT = 7'b0110011;
	parameter LD       = 7'b0000011;
	parameter SD       = 7'b0100011;
	parameter BEQ      = 7'b1100111;
	parameter ADDi     = 7'b0010011;
	parameter ORi      = 7'b0010011;

	always @(opcode) //when opcode is changed, following block is executed 
	begin
		case (opcode)
		// fill in the misisng code
		7'b0110011: begin
			ALUSrc <= 1'b0;
			MemtoReg <= 1'b0;
			RegWrite <= 1'b1;
			MemRead <= 1'b0;
			MemWrite <= 1'b0;
			Branch <= 1'b0;
			ALUOp <= 2'b10;
			end
		7'b0000011: begin
			ALUSrc <= 1'b1;
			MemtoReg <= 1'b1;
			RegWrite <= 1'b1;
			MemRead <= 1'b1;
			MemWrite <= 1'b0;
			Branch <= 1'b0;
			ALUOp <= 2'b00;
			end
		7'b0100011: begin
			ALUSrc <= 1'b1;
			MemtoReg <= 1'bx;
			RegWrite <= 1'b0;
			MemRead <= 1'b1;
			MemWrite <= 1'b1;
			Branch <= 1'b0;
			ALUOp <= 2'b00;
			end
		7'b1100111: begin
			ALUSrc <= 1'b0;
			MemtoReg <= 1'bx;
			RegWrite <= 1'b0;
			MemRead <= 1'b0;
			MemWrite <= 1'b0;
			Branch <= 1'b1;
			ALUOp <= 2'b01;
			end	
		7'b0010011: begin
			ALUSrc <= 1'b1;
			MemtoReg <= 1'b0;
			RegWrite <= 1'b1;
			MemRead <= 1'b0;
			MemWrite <= 1'b0;
			Branch <= 1'b0;
			ALUOp <= 2'b11;
			end
		// fill in the missing code  

		endcase
	end
endmodule

