library verilog;
use verilog.vl_types.all;
entity pr1_vlg_check_tst is
    port(
        X               : in     vl_logic;
        sampler_rx      : in     vl_logic
    );
end pr1_vlg_check_tst;
